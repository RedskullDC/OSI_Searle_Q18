
module first_nios1_system (
	clk_clk,
	reset_reset_n,
	pio_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pio_external_connection_export;
endmodule
